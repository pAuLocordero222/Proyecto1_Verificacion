class Envi #();
    

endclass